module LCD (input  Clk,
				input reset,
				output reg  [10:0]n_LCD_DATA,
				input [1:0]game_state
				);
reg  [10:0]LCD_DATA;	
reg [30:0]count;
reg [5:0]state;
reg [7:0]data[32:0];
always@ (posedge Clk or negedge reset) 
	begin
	if(~reset)
		begin
		count=30'd0;
		state=6'd0;
		n_LCD_DATA=11'b0;
		end
	else 
	begin
		if(game_state==1)state=0;
		if(game_state==2)state=0;
		if(count==25000)
			begin
			n_LCD_DATA=11'b0;
			if(state<40)state=state+1;
			count=0;
			LCD_DATA=11'b0;
			end
		else count=count+1;
		end
		n_LCD_DATA=LCD_DATA;
		case(state)
			6'd0:LCD_DATA=11'b00000000000;
			6'd1:LCD_DATA=11'b10000111000;
			6'd2:LCD_DATA=11'b10000001110;
			6'd3:LCD_DATA=11'b10000000001;
			6'd5:LCD_DATA=11'b10000000110;
			6'd6:LCD_DATA=11'b10010000000;
			6'd7:LCD_DATA={3'b110,data[0]};
			6'd8:LCD_DATA={3'b110,data[1]};
			6'd9:LCD_DATA={3'b110,data[2]};
			6'd10:LCD_DATA={3'b110,data[3]};
			6'd11:LCD_DATA={3'b110,data[4]};
			6'd12:LCD_DATA={3'b110,data[5]};
			6'd13:LCD_DATA={3'b110,data[6]};
			6'd14:LCD_DATA={3'b110,data[7]};
			6'd15:LCD_DATA={3'b110,data[8]};
			6'd16:LCD_DATA={3'b110,data[9]};
			6'd17:LCD_DATA={3'b110,data[10]};
			6'd18:LCD_DATA={3'b110,data[11]};
			6'd19:LCD_DATA={3'b110,data[12]};
			6'd20:LCD_DATA={3'b110,data[13]};
			6'd21:LCD_DATA={3'b110,data[14]};
			6'd22:LCD_DATA={3'b110,data[15]};
			6'd23:LCD_DATA=11'b10011000000;
			6'd24:LCD_DATA={3'b110,data[16]};
			6'd25:LCD_DATA={3'b110,data[17]};
			6'd26:LCD_DATA={3'b110,data[18]};
			6'd27:LCD_DATA={3'b110,data[19]};
			6'd28:LCD_DATA={3'b110,data[20]};
			6'd29:LCD_DATA={3'b110,data[21]};
			6'd30:LCD_DATA={3'b110,data[22]};
			6'd31:LCD_DATA={3'b110,data[23]};
			6'd32:LCD_DATA={3'b110,data[24]};
			6'd33:LCD_DATA={3'b110,data[25]};
			6'd34:LCD_DATA={3'b110,data[26]};
			6'd35:LCD_DATA={3'b110,data[27]};
			6'd36:LCD_DATA={3'b110,data[28]};
			6'd37:LCD_DATA={3'b110,data[29]};
			6'd38:LCD_DATA={3'b110,data[30]};
			6'd39:LCD_DATA={3'b110,data[31]};	
			default:LCD_DATA=11'b0;
		endcase
	end
always@ (game_state)begin
 if(game_state==0)begin
	  data[0]=8'b00100000;
	  data[1]=8'b01010000;//p
	  data[2]=8'b01101001;//i
	  data[3]=8'b01101110;//n
	  data[4]=8'b01100111;//g
	  data[5]=8'b00100000;
	  data[6]=8'b01010000;//p
	  data[7]=8'b01101111;//o
	  data[8]=8'b01101110;//n
	  data[9]=8'b01100111;//g
	  data[10]=8'b00100000;
	  data[11]=8'b00100000;
	  data[12]=8'b00100000;
	  data[13]=8'b00100000;
	  data[14]=8'b00100000;
	  data[15]=8'b00100000;
	  //
	  data[16]=8'b00100000;
	  data[17]=8'b00100000;
	  data[18]=8'b01000111;//G
	  data[19]=8'b01100001;//a
	  data[20]=8'b01101101;//m
	  data[21]=8'b01100101;//e
	  data[22]=8'b00100000;
	  data[23]=8'b00100000;
	  data[24]=8'b00100000;
	  data[25]=8'b00100000;
	  data[26]=8'b00100000;
	  data[27]=8'b00100000;
	  data[28]=8'b00100000;
	  data[29]=8'b00100000;
	  data[30]=8'b00100000;
	  data[31]=8'b00100000;
		end
 else if(game_state==1)begin
	  data[0]=8'b00100000;
	  data[1]=8'b01010000;//P
	  data[2]=8'b01101100;//l
	  data[3]=8'b01100001;//a
	  data[4]=8'b01111001;//y
	  data[5]=8'b01100101;//e
	  data[6]=8'b01110010;//r
	  data[7]=8'b00100000;// 
	  data[8]=8'b00100000;//
	  data[9]=8'b01000001;//A
	  data[10]=8'b00100000;
	  data[11]=8'b00100000;
	  data[12]=8'b00100000;
	  data[13]=8'b00100000;
	  data[14]=8'b00100000;
	  data[15]=8'b00100000;
	  //
	  data[16]=8'b00100000;
	  data[17]=8'b00100000;
	  data[18]=8'b01001001;//I
	  data[19]=8'b01110011;//s
	  data[20]=8'b00100000;//
	  data[21]=8'b01010111;//W
	  data[22]=8'b01101001;//i
	  data[23]=8'b01101110;//n
	  data[24]=8'b01101110;//n
	  data[25]=8'b01100101;//e
	  data[26]=8'b01110010;//r
	  data[27]=8'b00100001;//!
	  data[28]=8'b00100000;
	  data[29]=8'b00100000;
	  data[30]=8'b00100000;
	  data[31]=8'b00100000;
		end
 else if(game_state==2)begin
	  data[0]=8'b00100000;
	  data[1]=8'b01010000;//P
	  data[2]=8'b01101100;//l
	  data[3]=8'b01100001;//a
	  data[4]=8'b01111001;//y
	  data[5]=8'b01100101;//e
	  data[6]=8'b01110010;//r
	  data[7]=8'b00100000;// 
	  data[8]=8'b00100000;//
	  data[9]=8'b01000010;//B
	  data[10]=8'b00100000;
	  data[11]=8'b00100000;
	  data[12]=8'b00100000;
	  data[13]=8'b00100000;
	  data[14]=8'b00100000;
	  data[15]=8'b00100000;
	  //
	  data[16]=8'b00100000;
	  data[17]=8'b00100000;
	  data[18]=8'b01001001;//I
	  data[19]=8'b01110011;//s
	  data[20]=8'b00100000;//
	  data[21]=8'b01010111;//W
	  data[22]=8'b01101001;//i
	  data[23]=8'b01101110;//n
	  data[24]=8'b01101110;//n
	  data[25]=8'b01100101;//e
	  data[26]=8'b01110010;//r
	  data[27]=8'b00100001;//!
	  data[28]=8'b00100000;
	  data[29]=8'b00100000;
	  data[30]=8'b00100000;
	  data[31]=8'b00100000;
	end
end
endmodule
